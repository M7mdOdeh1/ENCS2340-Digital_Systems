//Name : Mohammed Owda
//id : 1200089
// BCD Adder using data flow

module BCD_Adder(a,b,cin,sum,cout)
input [3:0] a,b;
input cin,temp;